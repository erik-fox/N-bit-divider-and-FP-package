module top();

import 

endmodule
