module top();
import floatingpoint::*;

endmodule
